--Overflow
--verifica se a saida co da alu é 1 e da sinal pro controlador