--DataPath
--converter o RF_W_data de 8 pra 16 bits